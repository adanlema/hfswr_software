module bram_sincedge (
    input  wire     clk,
    input  wire     sinc,
    output wire     sinc_edge
);

//////////////////////////////////////////////////////////////////////////////////
//      WIRE AND REGISTERS
//////////////////////////////////////////////////////////////////////////////////
reg     sinc_prev;
reg     sinc_reg;

//////////////////////////////////////////////////////////////////////////////////
//      LOGICA
//////////////////////////////////////////////////////////////////////////////////
always @(posedge clk) begin
    // Almacenamos el valor previo de sinc
    sinc_prev <= sinc;
    
    // Comprobamos si hay un flanco ascendente en sinc
    if (sinc && !sinc_prev)
        sinc_reg <= 1'b1;
    else
        sinc_reg <= 1'b0;
end

//////////////////////////////////////////////////////////////////////////////////
//      SALIDAS
//////////////////////////////////////////////////////////////////////////////////
assign  sinc_edge   = sinc_reg;

endmodule
